library verilog;
use verilog.vl_types.all;
entity booth_alu_vlg_vec_tst is
end booth_alu_vlg_vec_tst;
