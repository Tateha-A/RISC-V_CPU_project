library ieee;
use ieee.std_logic_1164.all;

entity addi_tb is -- addi R2, R1, -5
end;